`timescale 1ns/1ps

module fibonacci_tb (clk, rst_n, en, sum);




endmodule 